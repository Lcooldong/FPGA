module tb_comb_gate;
    reg a, b, c, d, e;
    wire y;


    