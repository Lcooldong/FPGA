module and_gate(in1, in2, out1);
	
	input in1, in2;
	output out1;
	
	and(out1, in1, in2);
	
endmodule