module tb_dff;
    